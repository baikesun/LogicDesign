//	==================================================
//	Copyright (c) 2019 Sookmyung Women's University.
//	--------------------------------------------------
//	FILE 			: Project.v
//	DEPARTMENT		: EE
//	AUTHOR			: BAIK ESUN
//	EMAIL			: baik0705@sookmyung.ac.kr
//	--------------------------------------------------
//	RELEASE HISTORY
//	--------------------------------------------------
//	VERSION			DATE
//	0.0			2019-11-21
//	--------------------------------------------------
//	PURPOSE			: Digital Clock
//	==================================================

//	--------------------------------------------------
//	Numerical Controlled Oscillator
//	Hz of o_gen_clk = Clock Hz / num
//	--------------------------------------------------

module	nco(	
		o_gen_clk,
		i_nco_num,
		clk,
		rst_n);

	output		o_gen_clk	;	// 1Hz CLK

	input	[31:0]	i_nco_num	;
	input		clk		;	// 50Mhz CLK
	input		rst_n		;

	reg	[31:0]	cnt		;
	reg		o_gen_clk	;

	always @(posedge clk or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			cnt		<= 32'd0;
			o_gen_clk	<= 1'd0	;
		end 
		else begin
			if(cnt >= i_nco_num/2-1) begin
				cnt 	<= 32'd0		;
				o_gen_clk	<= ~o_gen_clk	;
			end 
			else begin
				cnt <= cnt + 1'b1		;
			end
		end
	end

endmodule

module	nco_down(	
		o_gen_clk,
		i_nco_num,
		clk,
		rst_n);

	output		o_gen_clk	;	// 1Hz CLK

	input	[31:0]	i_nco_num	;
	input		clk		;	// 50Mhz CLK
	input		rst_n		;

	reg	[31:0]	cnt		;
	reg		o_gen_clk	;

	always @(posedge clk or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			cnt		<= 32'd0;
			o_gen_clk	<= 1'd0	;
		end 
		else begin
			if(cnt <= 32'd0) begin
				cnt <= i_nco_num/2-1	;
				o_gen_clk <= ~o_gen_clk	;
			end 
			else begin
				cnt <= cnt - 1'b1	;
			end
		end
	end

endmodule

//	--------------------------------------------------
//	Flexible Numerical Display Decoder
//	--------------------------------------------------
module	fnd_dec(
		o_seg,
		i_num);

	output	[6:0]	o_seg		;	// {o_seg_a, o_seg_b, ... , o_seg_g}

	input	[3:0]	i_num		;

	reg	[6:0]	o_seg		;

	//making
	always @(i_num) begin 
	 	case(i_num) 
	 		4'd0 : o_seg = 7'b111_1110	; 
	 		4'd1 : o_seg = 7'b011_0000	; 
	 		4'd2 : o_seg = 7'b110_1101	; 
	 		4'd3 : o_seg = 7'b111_1001	; 
	 		4'd4 : o_seg = 7'b011_0011	; 
	 		4'd5 : o_seg = 7'b101_1011	; 
	 		4'd6 : o_seg = 7'b101_1111	; 
	 		4'd7 : o_seg = 7'b111_0000	; 
	 		4'd8 : o_seg = 7'b111_1111	; 
	 		4'd9 : o_seg = 7'b111_0011	; 
			default : o_seg = 7'b000_0000	; 
		endcase 
	end


endmodule

//	--------------------------------------------------
//	0~59 --> 2 Separated Segments
//	--------------------------------------------------
module	double_fig_sep(
		o_left,
		o_right,
		i_double_fig);

	output	[3:0]	o_left		;
	output	[3:0]	o_right		;
	
	input	[5:0]	i_double_fig	;
	
	assign		o_left	= i_double_fig / 10	;
	assign		o_right	= i_double_fig % 10	;
	
endmodule

//	--------------------------------------------------
//	0~59 --> 2 Separated Segments
//	--------------------------------------------------
module	led_disp(
		o_seg,
		o_seg_dp,
		o_seg_enb,
		i_six_digit_seg,
		i_six_dp,
		i_mode,
		i_position,
		clk,
		rst_n);

	output	[5:0]	o_seg_enb		;
	output		o_seg_dp		;
	output	[6:0]	o_seg			;
	
	input	[41:0]	i_six_digit_seg		;
	input	[5:0]	i_six_dp		;
	input	[2:0]	i_mode			;
	input	[1:0]	i_position		;

	input		clk			;
	input		rst_n			;

	parameter	MODE_CLOCK	= 3'd0	;
	parameter	MODE_SETUP	= 3'd1	;
	parameter	MODE_ALARM	= 3'd2	;
	parameter	MODE_TIMER_SET	= 3'd3	;
	parameter	MODE_TIMER	= 3'd4	;
	
	parameter	POS_SEC	= 2'd0		;
	parameter	POS_MIN	= 2'd1		;
	parameter	POS_HOU = 2'd2		;
	
	wire		gen_clk			;
	
	nco		u_nco(
			.o_gen_clk	(	gen_clk		),
			.i_nco_num	(	32'd5000	),
			.clk		(	clk		),
			.rst_n		(	rst_n		));

	wire		blink			;
	
	nco		u_nco_blink(
			.o_gen_clk	(	blink		),
			.i_nco_num	(	32'd100000000	),
			.clk		(	clk		),
			.rst_n		(	rst_n		));

	reg	[3:0]	cnt_common_node	;

	always @(posedge gen_clk or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			cnt_common_node <= 4'd0;
		end 
		else begin
			if(cnt_common_node >= 4'd5) begin
				cnt_common_node <= 4'd0;
			end 
			else begin
				cnt_common_node <= cnt_common_node + 1'b1;
			end
		end
	end
	
	reg	[5:0]	o_seg_enb		;

	always @(*) begin
		if ( (i_mode == MODE_SETUP) || (i_mode == MODE_ALARM) || (i_mode == MODE_TIMER_SET) ) begin
			case (i_position)
				POS_SEC : begin
					if ( blink == 1'b0 ) begin
						case (cnt_common_node)
							4'd0 	: o_seg_enb = 6'b111110;
							4'd1 	: o_seg_enb = 6'b111101;
							4'd2 	: o_seg_enb = 6'b111011;
							4'd3 	: o_seg_enb = 6'b110111;
							4'd4 	: o_seg_enb = 6'b101111;
							4'd5 	: o_seg_enb = 6'b011111;
							default	: o_seg_enb = 6'b111111;
						endcase
					end
					else begin
						case (cnt_common_node)
							4'd0 	: o_seg_enb = 6'b111111;
							4'd1 	: o_seg_enb = 6'b111111;
							4'd2 	: o_seg_enb = 6'b111011;
							4'd3 	: o_seg_enb = 6'b110111;
							4'd4 	: o_seg_enb = 6'b101111;
							4'd5 	: o_seg_enb = 6'b011111;
							default	: o_seg_enb = 6'b111111;
						endcase
					end
				end
				POS_MIN : begin
					if ( blink == 1'b0 ) begin
						case (cnt_common_node)
							4'd0 	: o_seg_enb = 6'b111110;
							4'd1 	: o_seg_enb = 6'b111101;
							4'd2 	: o_seg_enb = 6'b111011;
							4'd3 	: o_seg_enb = 6'b110111;
							4'd4 	: o_seg_enb = 6'b101111;
							4'd5 	: o_seg_enb = 6'b011111;
							default	: o_seg_enb = 6'b111111;
						endcase
					end
					else begin
						case (cnt_common_node)
							4'd0 	: o_seg_enb = 6'b111110;
							4'd1 	: o_seg_enb = 6'b111101;
							4'd2 	: o_seg_enb = 6'b111111;
							4'd3 	: o_seg_enb = 6'b111111;
							4'd4 	: o_seg_enb = 6'b101111;
							4'd5 	: o_seg_enb = 6'b011111;
							default	: o_seg_enb = 6'b111111;
						endcase
					end
				end
				POS_HOU : begin
					if ( blink == 1'b0 ) begin
						case (cnt_common_node)
							4'd0 	: o_seg_enb = 6'b111110;
							4'd1 	: o_seg_enb = 6'b111101;
							4'd2 	: o_seg_enb = 6'b111011;
							4'd3 	: o_seg_enb = 6'b110111;
							4'd4 	: o_seg_enb = 6'b101111;
							4'd5 	: o_seg_enb = 6'b011111;
							default	: o_seg_enb = 6'b111111;
						endcase
					end
					else begin
						case (cnt_common_node)
							4'd0 	: o_seg_enb = 6'b111110;
							4'd1 	: o_seg_enb = 6'b111101;
							4'd2 	: o_seg_enb = 6'b111011;
							4'd3 	: o_seg_enb = 6'b110111;
							4'd4 	: o_seg_enb = 6'b111111;
							4'd5 	: o_seg_enb = 6'b111111;
							default	: o_seg_enb = 6'b111111;
						endcase
					end
				end
			endcase
		end
		else begin
			case (cnt_common_node)
				4'd0 	: o_seg_enb = 6'b111110;
				4'd1 	: o_seg_enb = 6'b111101;
				4'd2 	: o_seg_enb = 6'b111011;
				4'd3 	: o_seg_enb = 6'b110111;
				4'd4 	: o_seg_enb = 6'b101111;
				4'd5 	: o_seg_enb = 6'b011111;
				default	: o_seg_enb = 6'b111111;
			endcase
		end
	end

	/*reg	[5:0]	o_seg_enb		;
	
	always @(cnt_common_node) begin
		case (cnt_common_node)
			4'd0 	: o_seg_enb = 6'b111110;
			4'd1 	: o_seg_enb = 6'b111101;
			4'd2 	: o_seg_enb = 6'b111011;
			4'd3 	: o_seg_enb = 6'b110111;
			4'd4 	: o_seg_enb = 6'b101111;
			4'd5 	: o_seg_enb = 6'b011111;
			default	: o_seg_enb = 6'b111111;
		endcase
	end*/
	
	reg		o_seg_dp		;

	always @(cnt_common_node) begin
		case (cnt_common_node)
			4'd0 	: o_seg_dp = i_six_dp[0];
			4'd1 	: o_seg_dp = i_six_dp[1];
			4'd2 	: o_seg_dp = i_six_dp[2];
			4'd3 	: o_seg_dp = i_six_dp[3];
			4'd4 	: o_seg_dp = i_six_dp[4];
			4'd5 	: o_seg_dp = i_six_dp[5];
			default	: o_seg_dp = 1'b0	;
		endcase
	end
	
	reg	[6:0]	o_seg			;

	always @(cnt_common_node) begin
		case (cnt_common_node)
			4'd0 	: o_seg = i_six_digit_seg[6:0]	;
			4'd1 	: o_seg = i_six_digit_seg[13:7]	;
			4'd2 	: o_seg = i_six_digit_seg[20:14];
			4'd3 	: o_seg = i_six_digit_seg[27:21];
			4'd4 	: o_seg = i_six_digit_seg[34:28];
			4'd5 	: o_seg = i_six_digit_seg[41:35];
			default	: o_seg = 7'b111_1110		;
		endcase
	end

endmodule

//	--------------------------------------------------
//	HMS(Hour:Min:Sec) Counter
//	--------------------------------------------------
module	hms_cnt(
		o_hms_cnt,
		o_max_hit,
		i_max_cnt,
		clk,
		rst_n);

	output	[5:0]	o_hms_cnt		;
	output		o_max_hit		;

	input	[5:0]	i_max_cnt		;
	input		clk			;
	input		rst_n			;

	reg	[5:0]	o_hms_cnt		;
	reg		o_max_hit		;

	always @(posedge clk or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			o_hms_cnt <= 6'd0;
			o_max_hit <= 1'b0;
		end 
		else begin
			if(o_hms_cnt >= i_max_cnt) begin
				o_hms_cnt <= 6'd0;
				o_max_hit <= 1'b1;
			end 
			else begin
				o_hms_cnt <= o_hms_cnt + 1'b1;
				o_max_hit <= 1'b0;
			end
		end
	end
endmodule

module	hms_cnt_down(
		o_hms_cnt,
		o_max_hit,
		i_max_cnt,
		clk,
		rst_n);

	output	[5:0]	o_hms_cnt		;
	output		o_max_hit		;

	input	[5:0]	i_max_cnt		;
	input		clk			;
	input		rst_n			;

	reg	[5:0]	o_hms_cnt		;
	reg		o_max_hit		;

	always @(posedge clk or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			o_hms_cnt <= 6'd0;
			o_max_hit <= 1'b0;
		end 
		else begin
			if(o_hms_cnt <= 6'd0) begin
				o_hms_cnt <= i_max_cnt;
				o_max_hit <= 1'b1;
			end 
			else begin
				o_hms_cnt <= o_hms_cnt - 1'b1;
				o_max_hit <= 1'b0;
			end
		end
	end

endmodule

module  debounce(
		o_sw,
		i_sw,
		clk);
	output		o_sw			;

	input		i_sw			;
	input		clk			;

	reg		dly1_sw			;

	always @(posedge clk) begin
		dly1_sw <= i_sw;
	end
	
	reg		dly2_sw			;

	always @(posedge clk) begin
		dly2_sw <= dly1_sw;
	end
	
	assign		o_sw = dly1_sw | ~dly2_sw;

endmodule

//	--------------------------------------------------
//	Clock Controller
//	--------------------------------------------------
module	controller(
		o_mode,
		o_position,
		o_alarm_en,
		o_timer_en,
		o_sec_clk,
		o_min_clk,
		o_hou_clk,
		o_alarm_sec_clk,
		o_alarm_min_clk,
		o_alarm_hou_clk,
		o_timer_sec_clk,
		o_timer_min_clk,
		o_timer_hou_clk,
		i_max_hit_sec,
		i_max_hit_min,
		i_max_hit_hou,
		i_max_hit_ts,
		i_max_hit_tm,
		i_sw0,
		i_sw1,
		i_sw2,
		i_sw3,
		i_sw4,
		clk,
		rst_n);

	output	[2:0]	o_mode			;
	output	[1:0]	o_position		;

	output		o_alarm_en		;
	output		o_timer_en		;

	output		o_sec_clk		;
	output		o_min_clk		;
	output		o_hou_clk		;

	output		o_alarm_sec_clk		;
	output		o_alarm_min_clk		;
	output		o_alarm_hou_clk		;

	output		o_timer_sec_clk		;
	output		o_timer_min_clk		;
	output		o_timer_hou_clk		;

	input		i_max_hit_sec		;
	input		i_max_hit_min		;
	input		i_max_hit_hou		;
	input		i_max_hit_ts		;
	input		i_max_hit_tm		;
	
	input		i_sw0			;
	input		i_sw1			;
	input		i_sw2			;
	input		i_sw3			;
	input		i_sw4			;
	
	input		clk			;
	input		rst_n			;

	parameter	MODE_CLOCK	= 3'd0	;
	parameter	MODE_SETUP	= 3'd1	;
	parameter	MODE_ALARM	= 3'd2	;
	parameter	MODE_TIMER_SET	= 3'd3	;
	parameter	MODE_TIMER	= 3'd4	;
	
	parameter	POS_SEC	= 2'd0		;
	parameter	POS_MIN	= 2'd1		;
	parameter	POS_HOU = 2'd2		;
	
	wire		clk_100hz		;

	nco		u0_nco(
			.o_gen_clk	( clk_100hz	),
			.i_nco_num	( 32'd500000	),
			.clk		( clk		),
			.rst_n		( rst_n		));
	
	wire		sw0			;

	debounce	u0_debounce(
			.o_sw		( sw0		),
			.i_sw		( i_sw0		),
			.clk		( clk_100hz	));
	
	wire		sw1			;

	debounce	u1_debounce(
			.o_sw		( sw1		),
			.i_sw		( i_sw1		),
			.clk		( clk_100hz	));
	
	wire		sw2			;

	debounce	u2_debounce(
			.o_sw		( sw2		),
			.i_sw		( i_sw2		),
			.clk		( clk_100hz	));

	wire		sw3			;

	debounce	u3_debounce(
			.o_sw		( sw3		),
			.i_sw		( i_sw3		),
			.clk		( clk_100hz	));

	wire		sw4			;

	debounce	u4_debounce(
			.o_sw		( sw4		),
			.i_sw		( i_sw4		),
			.clk		( clk_100hz	));
	
	reg	[2:0]	o_mode			;

	always @(posedge sw0 or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			o_mode <= MODE_CLOCK;
		end 
		else begin
			if(o_mode >= MODE_TIMER) begin
				o_mode <= MODE_CLOCK;
			end
			else begin
				o_mode <= o_mode + 1'b1;
			end
		end
	end

	reg	[1:0]	o_position		;

	always @(posedge sw1 or negedge rst_n) begin		//edit to change position directly to 'second' after 'hour'.
		if(rst_n == 1'b0) begin
			o_position <= POS_SEC;
		end 
		else begin
			if(o_position >= POS_HOU) begin
				o_position <= POS_SEC		;
			end
			else begin
				o_position <= o_position + 1'b1	;
			end 
		end
	end
	
	reg		o_alarm_en		;

	always @(posedge sw3 or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			o_alarm_en <= 1'b0;
		end 
		else begin
			o_alarm_en <= o_alarm_en + 1'b1;
		end
	end

	reg		o_timer_en		;

	always @(posedge sw4 or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			o_timer_en <= 1'b0;
		end
		else begin
			o_timer_en <= o_timer_en + 1'b1;
		end
	end

	wire		clk_1hz			;

	nco		u1_nco(
			.o_gen_clk	( clk_1hz	),
			.i_nco_num	( 32'd50000000	),
			.clk		( clk		),
			.rst_n		( rst_n		));

	wire		clk_down		;

	nco		u2_nco(
			.o_gen_clk	( clk_down	),
			.i_nco_num	( 32'd50000000	),
			.clk		( clk		),
			.rst_n		( rst_n		));
	
	reg		o_sec_clk		;
	reg		o_min_clk		;
	reg		o_hou_clk		;

	reg		o_alarm_sec_clk		;
	reg		o_alarm_min_clk		;
	reg		o_alarm_hou_clk		;

	reg		o_timer_sec_clk		;
	reg		o_timer_min_clk		;
	reg		o_timer_hou_clk		;

	always @(*) begin
		case(o_mode)
			MODE_CLOCK : begin
				o_sec_clk = clk_1hz;
				o_min_clk = i_max_hit_sec;
				o_hou_clk = i_max_hit_min;
				o_alarm_sec_clk = 1'b0;
				o_alarm_min_clk = 1'b0;
				o_alarm_hou_clk = 1'b0;
				o_timer_sec_clk = 1'b0;
				o_timer_min_clk = 1'b0;
				o_timer_hou_clk = 1'b0;
			end
			MODE_SETUP : begin
				case(o_position)
					POS_SEC : begin
						o_sec_clk = ~sw2;
						o_min_clk = 1'b0;
						o_hou_clk = 1'b0;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = 1'b0;
					end
					POS_MIN : begin
						o_sec_clk = 1'b0;
						o_min_clk = ~sw2;
						o_hou_clk = 1'b0;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = 1'b0;
					end
					POS_HOU : begin
						o_sec_clk = 1'b0;
						o_min_clk = 1'b0;
						o_hou_clk = ~sw2;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = 1'b0;
					end
						
				endcase
			end
			MODE_ALARM : begin
				case(o_position)
					POS_SEC : begin
						o_sec_clk = clk_1hz;
						o_min_clk = i_max_hit_sec;
						o_hou_clk = i_max_hit_min;
						o_alarm_sec_clk = ~sw2;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = 1'b0;
					end
					POS_MIN : begin
						o_sec_clk = clk_1hz;
						o_min_clk = i_max_hit_sec;
						o_hou_clk = i_max_hit_min;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = ~sw2;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = 1'b0;
					end
					POS_HOU : begin
						o_sec_clk = clk_1hz;
						o_min_clk = i_max_hit_sec;
						o_hou_clk = i_max_hit_min;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = ~sw2;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = 1'b0;
					end
				endcase
			end
			MODE_TIMER : begin
				if(o_timer_en == 1'b0) begin
					o_sec_clk = 1'b0;
					o_min_clk = 1'b0;
					o_hou_clk = 1'b0;
					o_alarm_sec_clk = 1'b0;
					o_alarm_min_clk = 1'b0;
					o_alarm_hou_clk = 1'b0;
					o_timer_sec_clk = 1'b0;
					o_timer_min_clk = 1'b0;
					o_timer_hou_clk = 1'b0;
				end
				else begin
					o_sec_clk = clk_1hz;
					o_min_clk = i_max_hit_sec;
					o_hou_clk = i_max_hit_min;
					o_alarm_sec_clk = 1'b0;
					o_alarm_min_clk = 1'b0;
					o_alarm_hou_clk = 1'b0;
					o_timer_sec_clk = clk_down;
					o_timer_min_clk = i_max_hit_ts;
					o_timer_hou_clk = i_max_hit_tm;
				end
			end
			MODE_TIMER_SET : begin
				case(o_position)
					POS_SEC : begin
						o_sec_clk = clk_1hz;
						o_min_clk = i_max_hit_sec;
						o_hou_clk = i_max_hit_min;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = ~sw2;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = 1'b0;
					end
					POS_MIN : begin
						o_sec_clk = clk_1hz;
						o_min_clk = i_max_hit_sec;
						o_hou_clk = i_max_hit_min;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = ~sw2;
						o_timer_hou_clk = 1'b0;
					end
					POS_HOU : begin
						o_sec_clk = clk_1hz;
						o_min_clk = i_max_hit_sec;
						o_hou_clk = i_max_hit_min;
						o_alarm_sec_clk = 1'b0;
						o_alarm_min_clk = 1'b0;
						o_alarm_hou_clk = 1'b0;
						o_timer_sec_clk = 1'b0;
						o_timer_min_clk = 1'b0;
						o_timer_hou_clk = ~sw2;
					end
				endcase
			end
			default : begin
				o_sec_clk = 1'b0;
				o_min_clk = 1'b0;
				o_hou_clk = 1'b0;
				o_alarm_sec_clk = 1'b0;
				o_alarm_min_clk = 1'b0;
				o_alarm_hou_clk = 1'b0;
				o_timer_sec_clk = 1'b0;
				o_timer_min_clk = 1'b0;
				o_timer_hou_clk = 1'b0;
			end
		endcase
	end

endmodule

//	--------------------------------------------------
//	HMS(Hour:Min:Sec) Counter
//	--------------------------------------------------
module	minsec(	o_sec,
		o_min,
		o_hou,
		o_max_hit_sec,
		o_max_hit_min,
		o_max_hit_hou,
		o_max_hit_ts,
		o_max_hit_tm,
		o_alarm,
		o_timer,
		i_mode,
		i_position,
		i_sec_clk,
		i_min_clk,
		i_hou_clk,
		i_alarm_sec_clk,
		i_alarm_min_clk,
		i_alarm_hou_clk,
		i_timer_sec_clk,
		i_timer_min_clk,
		i_timer_hou_clk,
		i_alarm_en,
		i_timer_en,
		clk,
		rst_n);

	output	[5:0]	o_sec		;
	output	[5:0]	o_min		;
	output	[5:0]	o_hou		;
	output		o_max_hit_sec	;
	output		o_max_hit_min	;
	output		o_max_hit_hou	;
	output		o_max_hit_ts	;
	output		o_max_hit_tm	;
	output		o_alarm		;
	output		o_timer		;
	
	input	[2:0]	i_mode		;
	input		i_position	;
	input		i_sec_clk	;
	input		i_min_clk	;
	input		i_hou_clk	;
	input		i_alarm_sec_clk	;
	input		i_alarm_min_clk	;
	input		i_alarm_hou_clk	;
	input		i_timer_sec_clk	;
	input		i_timer_min_clk	;
	input		i_timer_hou_clk	;
	input		i_alarm_en	;
	input		i_timer_en	;
	
	input		clk		;
	input		rst_n		;

	parameter	MODE_CLOCK	= 3'd0	;
	parameter	MODE_SETUP	= 3'd1	;
	parameter	MODE_ALARM	= 3'd2	;
	parameter	MODE_TIMER_SET	= 3'd3	;
	parameter	MODE_TIMER	= 3'd4	;

	parameter	POS_SEC		= 2'b00	;
	parameter	POS_MIN		= 2'b01	;
	parameter	POS_HOU		= 2'b10	;

	//MODE_CLOCK
	wire	[5:0]	sec		;
	wire		o_max_hit_sec	;
	
	hms_cnt		u0_hms_cnt(
				.o_hms_cnt	(	sec		),
				.o_max_hit	(	o_max_hit_sec	),
				.i_max_cnt	(	6'd59		),
				.clk		(	i_sec_clk	),
				.rst_n		(	rst_n		));
	
	wire	[5:0]	min		;
	wire		o_max_hit_min	;

	hms_cnt		u1_hms_cnt(
				.o_hms_cnt	(	min		),
				.o_max_hit	(	o_max_hit_min	),
				.i_max_cnt	(	6'd59		),
				.clk		(	i_min_clk	),
				.rst_n		(	rst_n		));

	wire	[5:0]	hou		;
	wire		o_max_hit_hou	;

	hms_cnt		u2_hms_cnt(
				.o_hms_cnt	(	hou		),
				.o_max_hit	(	o_max_hit_hou	),
				.i_max_cnt	(	6'd23		),
				.clk		(	i_hou_clk	),
				.rst_n		(	rst_n		));

	

	//	MODE_ALARM
	wire	[5:0]	alarm_sec	;

	hms_cnt		u_hms_cnt_alarm_sec(
				.o_hms_cnt	(	alarm_sec	),
				.o_max_hit	( 			),
				.i_max_cnt	(	6'd59		),
				.clk		(	i_alarm_sec_clk	),
				.rst_n		(	rst_n		));

	wire	[5:0]	alarm_min	;

	hms_cnt		u_hms_cnt_alarm_min(
				.o_hms_cnt	(	alarm_min	),
				.o_max_hit	( 			),
				.i_max_cnt	(	6'd59		),
				.clk		(	i_alarm_min_clk	),
				.rst_n		(	rst_n		));
	
	wire	[5:0]	alarm_hou	;

	hms_cnt		u_hms_cnt_alarm_hou(
				.o_hms_cnt	(	alarm_hou	),
				.o_max_hit	( 			),
				.i_max_cnt	(	6'd23		),
				.clk		(	i_alarm_hou_clk	),
				.rst_n		(	rst_n		));

	//	MODE_TIMER
	wire	[5:0]	timer_sec	;
	wire		o_max_hit_ts	;

	hms_cnt_down	u_hms_cnt_timer_sec(
				.o_hms_cnt	(	timer_sec	),
				.o_max_hit	( 	o_max_hit_ts	),
				.i_max_cnt	(	6'd59		),
				.clk		(	i_timer_sec_clk	),
				.rst_n		(	rst_n		));

	wire	[5:0]	timer_min	;
	wire		o_max_hit_tm	;

	hms_cnt_down	u_hms_cnt_timer_min(
				.o_hms_cnt	(	timer_min	),
				.o_max_hit	( 	o_max_hit_tm	),
				.i_max_cnt	(	6'd59		),
				.clk		(	i_timer_min_clk	),
				.rst_n		(	rst_n		));
	
	wire	[5:0]	timer_hou	;

	hms_cnt_down	u_hms_cnt_timer_hou(
				.o_hms_cnt	(	timer_hou	),
				.o_max_hit	( 			),
				.i_max_cnt	(	6'd23		),
				.clk		(	i_timer_hou_clk	),
				.rst_n		(	rst_n		));

	reg	[5:0]	o_sec		;
	reg	[5:0]	o_min		;
	reg	[5:0]	o_hou		;

	always @ (*) begin
		case(i_mode)
			MODE_CLOCK: 	begin
				o_sec	= sec;
				o_min	= min;
				o_hou	= hou;
			end
			MODE_SETUP:	begin
				o_sec	= sec;
				o_min	= min;
				o_hou	= hou;
			end
			MODE_ALARM:	begin
				o_sec	= alarm_sec;
				o_min	= alarm_min;
				o_hou	= alarm_hou;
			end
			MODE_TIMER:	begin
				o_sec	= timer_sec;
				o_min	= timer_min;
				o_hou	= timer_hou;
			end
			MODE_TIMER_SET:	begin
				o_sec	= timer_sec;
				o_min	= timer_min;
				o_hou	= timer_hou;
			end
		endcase
	end

	reg		o_alarm		;

	always @ (posedge clk or negedge rst_n) begin
		if (rst_n == 1'b0) begin
			o_alarm <= 1'b0;
		end 
		else begin
			if( (sec == alarm_sec) && (min == alarm_min) && (hou == alarm_hou)) begin
				o_alarm <= 1'b1 & i_alarm_en;
			end 
			else begin
				o_alarm <= o_alarm & i_alarm_en;
			end
		end
	end

	reg		o_timer		;

	always @ (posedge clk or negedge rst_n) begin
		if (rst_n == 1'b0) begin
			o_timer <= 1'b0;
		end 
		else begin
			if( (timer_sec == 6'd0) && (timer_min == 6'd0) && (timer_hou == 6'd0)) begin
				o_timer <= 1'b1 & i_timer_en;
			end 
			else begin
				o_timer <= o_timer & i_timer_en;
			end
		end
	end
endmodule

module	buzz(
		o_buzz,
		i_buzz_en1,
		i_buzz_en2,
		clk,
		rst_n);

	output		o_buzz		;

	input		i_buzz_en1	;	//alarm enable
	input		i_buzz_en2	;	//timer enable
	input		clk		;
	input		rst_n		;

	parameter	C = 191113	;
	parameter	D = 170262	;
	parameter	E = 151686	;
	parameter	F = 143173	;
	parameter	G = 63776	;
	parameter	A = 56818	;
	parameter	B = 50619	;

	wire		clk_beat		;

	nco	u_nco_beat(	
			.o_gen_clk	(	clk_beat		),
			.i_nco_num	(	25000000	),	//2Hz
			.clk		(	clk		),
			.rst_n		(	rst_n		));

	reg	[4:0]	cnt		;

	always @ (posedge clk_beat or negedge rst_n) begin
		if(rst_n == 1'b0) begin
			cnt <= 5'd0;
		end
		else begin
			if( (i_buzz_en1 == 1'b0) && (i_buzz_en2 == 1'b0) ) begin
				cnt <= 5'b0;
			end
			else begin
				if(cnt >= 5'd24) begin
					cnt <= 5'd0;
				end
				else begin
					cnt <= cnt + 1'd1;
				end
			end
		end
	end

	reg	[31:0]	nco_num		;

	always @ (*) begin
		case(cnt)
			5'd00: nco_num = E	;
			5'd01: nco_num = D	;
			5'd02: nco_num = C	;
			5'd03: nco_num = D	;
			5'd04: nco_num = E	;
			5'd05: nco_num = E	;
			5'd06: nco_num = E	;
			5'd07: nco_num = D	;
			5'd08: nco_num = D	;
			5'd09: nco_num = D	;
			5'd10: nco_num = E	;
			5'd11: nco_num = E	;
			5'd12: nco_num = E	;
			5'd13: nco_num = E	;
			5'd14: nco_num = D	;
			5'd15: nco_num = C	;
			5'd16: nco_num = D	;
			5'd17: nco_num = E	;
			5'd18: nco_num = E	;
			5'd19: nco_num = E	;
			5'd20: nco_num = D	;
			5'd21: nco_num = D	;
			5'd22: nco_num = E	;
			5'd23: nco_num = D	;
			5'd24: nco_num = C	;
		endcase
	end

	wire		buzz		;
	nco	u_nco_buzz(	
			.o_gen_clk	(	buzz		),
			.i_nco_num	(	nco_num		),
			.clk		(	clk		),
			.rst_n		(	rst_n		));

	assign		o_buzz = buzz & ( i_buzz_en1 | i_buzz_en2 );

	endmodule

module	top(
		o_seg_enb,
		o_seg_dp,
		o_seg,
		o_alarm,
		i_sw0,
		i_sw1,
		i_sw2,
		i_sw3,
		i_sw4,
		clk,
		rst_n);

	output	[5:0]	o_seg_enb	;
	output		o_seg_dp	;
	output	[6:0]	o_seg		;
	output		o_alarm		;
	
	input		i_sw0		;
	input		i_sw1		;
	input		i_sw2		;
	input		i_sw3		;
	input		i_sw4		;
	input		clk		;
	input		rst_n		;

	wire	[2:0]	mode		;
	wire	[1:0]	position	;
	wire		alarm_enb	;
	wire		timer_enb	;
	wire		alarm_hou_clk	;
	wire		alarm_min_clk	;
	wire		alarm_sec_clk	;
	wire		max_hit_hou	;
	wire		max_hit_min	;
	wire		max_hit_sec	;
	wire		max_hit_ts	;
	wire		max_hit_tm	;
	wire		hou_clk		;
	wire		min_clk		;
	wire		sec_clk		;

	controller	u_ctrl		(
						.o_mode			(	mode		),
						.o_position		(	position	),
						.o_alarm_en		(	alarm_enb	),
						.o_timer_en		(	timer_enb	),
						.o_sec_clk		(	sec_clk		),
						.o_min_clk		(	min_clk		),
						.o_hou_clk		(	hou_clk		),
						.o_alarm_sec_clk	(	alarm_sec_clk	),
						.o_alarm_min_clk	(	alarm_min_clk	),
						.o_alarm_hou_clk	(	alarm_hou_clk	),
						.o_timer_sec_clk	(	timer_sec_clk	),
						.o_timer_min_clk	(	timer_min_clk	),
						.o_timer_hou_clk	(	timer_hou_clk	),
						.i_max_hit_sec		(	max_hit_sec	),
						.i_max_hit_min		(	max_hit_min	),
						.i_max_hit_hou		(	max_hit_hou	),
						.i_max_hit_ts		(	max_hit_ts	),
						.i_max_hit_tm		(	max_hit_tm	),
						.i_sw0			(	i_sw0		),
						.i_sw1			(	i_sw1		),
						.i_sw2			(	i_sw2		),
						.i_sw3			(	i_sw3		),
						.i_sw4			(	i_sw4		),
						.clk			(	clk		),
						.rst_n			(	rst_n		));

	wire	[5:0]	hou		;	
	wire	[5:0]	min		;
	wire	[5:0]	sec		;
	wire		alarm		;
	wire		timer		;

	minsec		u_minsec	(	
						.o_sec			(	sec		),
						.o_min			(	min		),
						.o_hou			(	hou		),
						.o_max_hit_sec		(	max_hit_sec	),
						.o_max_hit_min		(	max_hit_min	),
						.o_max_hit_hou		(	max_hit_hou	),
						.o_max_hit_ts		(	max_hit_ts	),
						.o_max_hit_tm		(	max_hit_tm	),
						.o_alarm		(	alarm		),
						.o_timer		(	timer		),
						.i_mode			(	mode		),
						.i_position		(	position	),
						.i_sec_clk		(	sec_clk		),
						.i_min_clk		(	min_clk		),
						.i_hou_clk		(	hou_clk		),
						.i_alarm_sec_clk	(	alarm_sec_clk	),
						.i_alarm_min_clk	(	alarm_min_clk	),
						.i_alarm_hou_clk	(	alarm_hou_clk	),
						.i_timer_sec_clk	(	timer_sec_clk	),
						.i_timer_min_clk	(	timer_min_clk	),
						.i_timer_hou_clk	(	timer_hou_clk	),
						.i_alarm_en		(	alarm_enb	),
						.i_timer_en		(	timer_enb	),
						.clk			(	clk		),
						.rst_n			(	rst_n		));

	wire	[3:0]	sec_left	;
	wire	[3:0]	sec_right	;

	double_fig_sep	u0_dfs		(
						.o_left			(	sec_left	),
						.o_right		(	sec_right	),
						.i_double_fig		(	sec		));

	wire	[3:0]	min_left	;
	wire	[3:0]	min_right	;

	double_fig_sep	u1_dfs		(
						.o_left			(	min_left	),
						.o_right		(	min_right	),
						.i_double_fig		(	min		));

	wire	[3:0]	hou_left	;
	wire	[3:0]	hou_right	;

	double_fig_sep	u2_dfs		(
						.o_left			(	hou_left	),
						.o_right		(	hou_right	),
						.i_double_fig		(	hou		));

	wire	[6:0]	seg_first	;   //sec_right
	wire	[6:0]	seg_second	;   //sec_left
	wire	[6:0]	seg_third	;   //min_right
	wire	[6:0]	seg_fourth	;   //min_left
	wire	[6:0]	seg_fifth	;   //hou_right
	wire	[6:0]	seg_sixth	;   //hou_left

	fnd_dec		u0_fnd_dec	(
						.o_seg			(	seg_second	),
						.i_num			(	sec_left	));

	fnd_dec		u1_fnd_dec	(
						.o_seg			(	seg_first	),
						.i_num			(	sec_right	));

	fnd_dec		u2_fnd_dec	(
						.o_seg			(	seg_fourth	),
						.i_num			(	min_left	));

	fnd_dec		u3_fnd_dec	(
						.o_seg			(	seg_third	),
						.i_num			(	min_right	));

	fnd_dec		u4_fnd_dec	(
						.o_seg			(	seg_sixth	),
						.i_num			(	hou_left	));

	fnd_dec		u5_fnd_dec	(
						.o_seg			(	seg_fifth	),
						.i_num			(	hou_right	));

	wire	[41:0]	six_digit_seg	;
	
	assign		six_digit_seg = {seg_sixth, seg_fifth, seg_fourth, seg_third, seg_second, seg_first}	;

	led_disp	u_led_disp	(
						.o_seg			(	o_seg		),
						.o_seg_dp		(	o_seg_dp	),
						.o_seg_enb		(	o_seg_enb	),
						.i_six_digit_seg	(	six_digit_seg	),
						.i_six_dp		(	mode		),
						.i_mode			(	mode		),
						.i_position		(	position	),
						.clk			(	clk		),
						.rst_n			(	rst_n		));

	buzz		u_buzz		(
						.o_buzz			(	o_alarm		),
						.i_buzz_en1		(	alarm		),
						.i_buzz_en2		(	timer		),
						.clk			(	clk		),
						.rst_n			(	rst_n		));
	
endmodule
